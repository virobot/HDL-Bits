module top_module(
    input clk,
    input [7:0] in,
    input reset,    // Synchronous reset
    output [23:0] out_bytes,
    output done); //
	parameter BYTE1=0,BYTE2=1,BYTE3=2,DONE=3;
    reg [1:0] state,next_state;
    reg [23:0] data;
    // FSM from fsm_ps2
    always @(*) begin
        case(state)
            BYTE1 : next_state = (in[3]) ? BYTE2: BYTE1;
            BYTE2 : next_state = BYTE3;
            BYTE3 : next_state = DONE;
            DONE : next_state = (in[3]) ? BYTE2 : BYTE1;
        endcase
    end
    
    always @(posedge clk) begin
        if(reset) begin
            state<=BYTE1;
        	data<=24'b0;
        end
        else begin
            state<=next_state;
            data<={data[15:8],data[7:0],in};
        end
    end
    
    // New: Datapath to store incoming bytes.
    assign done = (state == DONE);
    assign out_bytes = (DONE) ? data : 24'b0;
endmodule
