module top_module(input a,b,c, output x,y,w,z);
	assign w=a,x=b,y=b,z=c;
endmodule